magic
tech sky130A
magscale 1 2
timestamp 1729050412
<< error_s >>
rect 170 2156 176 2162
rect 302 2156 308 2162
rect 164 2150 170 2156
rect 308 2154 314 2156
rect 2532 2154 2538 2160
rect 2538 2148 2544 2154
rect 164 2088 170 2094
rect 170 2082 176 2088
rect 2406 2074 2412 2080
rect 2538 2074 2544 2080
rect 2412 2068 2418 2074
rect 2532 2068 2538 2074
<< viali >>
rect 328 2598 2512 2752
rect 302 1494 2470 1648
<< metal1 >>
rect 316 2752 2524 2758
rect 316 2598 328 2752
rect 2512 2598 2524 2752
rect 316 2592 2524 2598
rect 162 2156 320 2160
rect 162 2088 170 2156
rect 308 2088 320 2156
rect 2402 2154 2552 2164
rect 890 2096 1112 2140
rect 162 2080 320 2088
rect 1692 2080 1892 2152
rect 2402 2074 2412 2154
rect 2538 2074 2552 2154
rect 2402 2068 2552 2074
rect 290 1648 2482 1654
rect 290 1494 302 1648
rect 2470 1494 2482 1648
rect 290 1488 2482 1494
<< via1 >>
rect 170 2088 308 2156
rect 2412 2074 2538 2154
<< metal2 >>
rect 308 2088 2412 2154
rect 176 2086 2412 2088
use inverter  x1
timestamp 1728978927
transform 1 0 53 0 1 1306
box 232 246 866 1374
use inverter  x2
timestamp 1728978927
transform 1 0 844 0 1 1306
box 232 246 866 1374
use inverter  x3
timestamp 1728978927
transform 1 0 1635 0 1 1306
box 232 246 866 1374
<< labels >>
flabel viali 396 2718 396 2718 0 FreeSans 800 0 0 0 vdd
port 0 nsew
flabel viali 362 1546 380 1582 0 FreeSans 800 0 0 0 gnd
port 1 nsew
flabel via1 2470 2110 2522 2142 0 FreeSans 800 0 0 0 out
port 2 nsew
<< end >>
