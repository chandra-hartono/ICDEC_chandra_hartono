magic
tech sky130A
magscale 1 2
timestamp 1729219852
<< nmos >>
rect -229 109 -29 509
rect 29 109 229 509
rect -229 -509 -29 -109
rect 29 -509 229 -109
<< ndiff >>
rect -287 497 -229 509
rect -287 121 -275 497
rect -241 121 -229 497
rect -287 109 -229 121
rect -29 497 29 509
rect -29 121 -17 497
rect 17 121 29 497
rect -29 109 29 121
rect 229 497 287 509
rect 229 121 241 497
rect 275 121 287 497
rect 229 109 287 121
rect -287 -121 -229 -109
rect -287 -497 -275 -121
rect -241 -497 -229 -121
rect -287 -509 -229 -497
rect -29 -121 29 -109
rect -29 -497 -17 -121
rect 17 -497 29 -121
rect -29 -509 29 -497
rect 229 -121 287 -109
rect 229 -497 241 -121
rect 275 -497 287 -121
rect 229 -509 287 -497
<< ndiffc >>
rect -275 121 -241 497
rect -17 121 17 497
rect 241 121 275 497
rect -275 -497 -241 -121
rect -17 -497 17 -121
rect 241 -497 275 -121
<< poly >>
rect -229 581 -29 597
rect -229 547 -213 581
rect -45 547 -29 581
rect -229 509 -29 547
rect 29 581 229 597
rect 29 547 45 581
rect 213 547 229 581
rect 29 509 229 547
rect -229 71 -29 109
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 109
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -109 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -109 229 -71
rect -229 -547 -29 -509
rect -229 -581 -213 -547
rect -45 -581 -29 -547
rect -229 -597 -29 -581
rect 29 -547 229 -509
rect 29 -581 45 -547
rect 213 -581 229 -547
rect 29 -597 229 -581
<< polycont >>
rect -213 547 -45 581
rect 45 547 213 581
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -213 -581 -45 -547
rect 45 -581 213 -547
<< locali >>
rect -229 547 -213 581
rect -45 547 -29 581
rect 29 547 45 581
rect 213 547 229 581
rect -275 497 -241 513
rect -275 105 -241 121
rect -17 497 17 513
rect -17 105 17 121
rect 241 497 275 513
rect 241 105 275 121
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect -275 -121 -241 -105
rect -275 -513 -241 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 241 -121 275 -105
rect 241 -513 275 -497
rect -229 -581 -213 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 213 -581 229 -547
<< viali >>
rect -213 547 -45 581
rect 45 547 213 581
rect -275 121 -241 497
rect -17 121 17 497
rect 241 121 275 497
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -275 -497 -241 -121
rect -17 -497 17 -121
rect 241 -497 275 -121
rect -213 -581 -45 -547
rect 45 -581 213 -547
<< metal1 >>
rect -225 581 -33 587
rect -225 547 -213 581
rect -45 547 -33 581
rect -225 541 -33 547
rect 33 581 225 587
rect 33 547 45 581
rect 213 547 225 581
rect 33 541 225 547
rect -281 497 -235 509
rect -281 121 -275 497
rect -241 121 -235 497
rect -281 109 -235 121
rect -23 497 23 509
rect -23 121 -17 497
rect 17 121 23 497
rect -23 109 23 121
rect 235 497 281 509
rect 235 121 241 497
rect 275 121 281 497
rect 235 109 281 121
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect -281 -121 -235 -109
rect -281 -497 -275 -121
rect -241 -497 -235 -121
rect -281 -509 -235 -497
rect -23 -121 23 -109
rect -23 -497 -17 -121
rect 17 -497 23 -121
rect -23 -509 23 -497
rect 235 -121 281 -109
rect 235 -497 241 -121
rect 275 -497 281 -121
rect 235 -509 281 -497
rect -225 -547 -33 -541
rect -225 -581 -213 -547
rect -45 -581 -33 -547
rect -225 -587 -33 -581
rect 33 -547 225 -541
rect 33 -581 45 -547
rect 213 -581 225 -547
rect 33 -587 225 -581
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 2 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
