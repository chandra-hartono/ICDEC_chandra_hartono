magic
tech sky130A
magscale 1 2
timestamp 1729397135
<< nwell >>
rect -176 -694 1280 562
<< nsubdiff >>
rect -140 492 -83 526
rect 1184 492 1244 526
rect -140 466 -106 492
rect 1210 466 1244 492
rect -140 -624 -106 -598
rect 1210 -624 1244 -598
rect -140 -658 -83 -624
rect 1184 -658 1244 -624
<< nsubdiffcont >>
rect -83 492 1184 526
rect -140 -598 -106 466
rect 1210 -598 1244 466
rect -83 -658 1184 -624
<< poly >>
rect -56 400 10 401
rect -56 385 37 400
rect -56 351 -40 385
rect -6 351 37 385
rect 1067 384 1154 400
rect -56 326 37 351
rect 382 346 721 380
rect 1067 350 1107 384
rect 1141 350 1154 384
rect 1067 325 1154 350
rect -79 -480 35 -447
rect -79 -493 -45 -480
rect -78 -514 -45 -493
rect -11 -514 35 -480
rect 382 -509 722 -475
rect 1068 -476 1155 -450
rect -78 -534 35 -514
rect 1068 -510 1105 -476
rect 1139 -510 1155 -476
rect 1068 -521 1155 -510
rect 1099 -523 1155 -521
<< polycont >>
rect -40 351 -6 385
rect 1107 350 1141 384
rect -45 -514 -11 -480
rect 1105 -510 1139 -476
<< locali >>
rect -140 492 -83 526
rect 1184 492 1244 526
rect -140 466 -106 492
rect 1210 466 1244 492
rect -56 351 -40 385
rect -6 351 10 385
rect 1095 384 1156 400
rect -49 314 6 351
rect 1091 350 1107 384
rect 1141 350 1156 384
rect -51 247 6 314
rect 1095 246 1156 350
rect -49 -370 9 -367
rect -49 -480 10 -370
rect 1100 -468 1148 -402
rect -51 -514 -45 -480
rect -11 -514 10 -480
rect -49 -533 10 -514
rect 1084 -476 1148 -468
rect 1084 -510 1105 -476
rect 1139 -510 1155 -476
rect 1084 -512 1148 -510
rect 1084 -521 1144 -512
rect -140 -624 -106 -598
rect 1210 -624 1244 -598
rect -140 -658 -83 -624
rect 1184 -658 1244 -624
<< viali >>
rect -40 351 -6 385
rect 1107 350 1141 384
rect 1206 -126 1210 -78
rect 1210 -126 1244 -78
rect 1244 -126 1250 -78
rect -45 -514 -11 -480
rect 1105 -510 1139 -476
<< metal1 >>
rect 126 454 671 455
rect 126 422 976 454
rect -52 385 6 391
rect -52 351 -40 385
rect -6 351 6 385
rect 126 381 159 422
rect -52 345 6 351
rect -49 314 6 345
rect 105 327 115 381
rect 173 327 183 381
rect 652 329 662 381
rect 714 329 724 381
rect 944 347 976 422
rect 1095 384 1156 400
rect 1095 350 1107 384
rect 1141 350 1156 384
rect -51 298 6 314
rect 1095 302 1156 350
rect -51 247 82 298
rect -48 157 82 247
rect -48 108 41 157
rect 31 98 41 108
rect 106 98 116 157
rect 205 111 351 287
rect 475 172 627 294
rect 475 120 527 172
rect 579 120 627 172
rect 227 -242 338 111
rect 475 104 627 120
rect 751 112 898 288
rect 1020 246 1156 302
rect 1020 161 1142 246
rect 767 -241 882 112
rect 1003 107 1013 161
rect 1065 108 1142 161
rect 1065 107 1075 108
rect 1200 -78 1256 -66
rect 1200 -126 1206 -78
rect 1250 -126 1256 -78
rect 1200 -138 1256 -126
rect -42 -254 84 -242
rect -42 -310 38 -254
rect 90 -310 100 -254
rect -42 -367 84 -310
rect -49 -420 84 -367
rect 206 -328 352 -242
rect 206 -380 254 -328
rect 306 -380 352 -328
rect 206 -418 352 -380
rect 480 -296 627 -243
rect 480 -352 519 -296
rect 581 -352 627 -296
rect 480 -419 627 -352
rect 750 -326 897 -241
rect 1014 -273 1140 -240
rect 1001 -325 1011 -273
rect 1063 -325 1140 -273
rect 750 -390 788 -326
rect 858 -390 897 -326
rect 750 -419 897 -390
rect 1014 -402 1140 -325
rect 1014 -418 1148 -402
rect -49 -474 10 -420
rect -51 -480 10 -474
rect -51 -514 -45 -480
rect -11 -514 10 -480
rect -51 -520 10 -514
rect -49 -533 10 -520
rect 128 -546 161 -476
rect 380 -510 390 -458
rect 442 -510 452 -458
rect 925 -510 935 -458
rect 987 -510 997 -458
rect 1100 -468 1148 -418
rect 1084 -470 1148 -468
rect 1084 -476 1151 -470
rect 1084 -510 1105 -476
rect 1139 -510 1151 -476
rect 945 -546 978 -510
rect 1084 -516 1151 -510
rect 1084 -521 1144 -516
rect 128 -579 978 -546
<< via1 >>
rect 115 327 173 381
rect 662 329 714 381
rect 41 98 106 157
rect 527 120 579 172
rect 1013 107 1065 161
rect 38 -310 90 -254
rect 254 -380 306 -328
rect 519 -352 581 -296
rect 1011 -325 1063 -273
rect 788 -390 858 -326
rect 390 -510 442 -458
rect 935 -510 987 -458
<< metal2 >>
rect -40 422 161 457
rect -40 -94 -5 422
rect 126 391 161 422
rect 662 454 714 455
rect 662 423 1144 454
rect 115 381 173 391
rect 115 317 173 327
rect 662 381 714 423
rect 662 319 714 329
rect 525 176 581 186
rect 41 157 106 167
rect 40 98 41 121
rect 525 110 581 120
rect 1013 161 1065 171
rect 40 88 106 98
rect 1013 97 1065 107
rect 40 -12 73 88
rect 519 -12 583 -10
rect 1021 -12 1054 97
rect 40 -45 1054 -12
rect 40 -49 73 -45
rect -38 -547 -5 -94
rect 38 -254 94 -244
rect 519 -296 583 -45
rect 1011 -269 1063 -263
rect 38 -320 94 -310
rect 224 -316 336 -306
rect 581 -352 583 -296
rect 519 -361 583 -352
rect 764 -314 876 -304
rect 1002 -325 1011 -269
rect 1067 -325 1076 -269
rect 519 -362 581 -361
rect 224 -404 336 -394
rect 1011 -335 1063 -325
rect 764 -402 876 -392
rect 390 -458 442 -448
rect 390 -516 442 -510
rect 935 -458 987 -448
rect 401 -547 434 -516
rect 935 -520 987 -510
rect -38 -580 434 -547
rect 937 -547 987 -520
rect 1109 -547 1140 423
rect 937 -578 1140 -547
rect 937 -579 987 -578
<< via2 >>
rect 525 172 581 176
rect 525 120 527 172
rect 527 120 579 172
rect 579 120 581 172
rect 38 -310 90 -254
rect 90 -310 94 -254
rect 224 -328 336 -316
rect 224 -380 254 -328
rect 254 -380 306 -328
rect 306 -380 336 -328
rect 764 -326 876 -314
rect 1011 -273 1067 -269
rect 1011 -325 1063 -273
rect 1063 -325 1067 -273
rect 224 -394 336 -380
rect 764 -390 788 -326
rect 788 -390 858 -326
rect 858 -390 876 -326
rect 764 -392 876 -390
<< metal3 >>
rect 515 176 591 181
rect 515 120 525 176
rect 581 120 591 176
rect 515 115 591 120
rect 518 -56 590 115
rect 10 -120 1071 -56
rect 10 -190 74 -120
rect 10 -194 105 -190
rect 9 -254 105 -194
rect 9 -310 38 -254
rect 94 -310 105 -254
rect 1007 -264 1071 -120
rect 1006 -269 1072 -264
rect 9 -325 105 -310
rect 214 -316 346 -311
rect 214 -394 224 -316
rect 336 -394 346 -316
rect 214 -399 346 -394
rect 754 -314 886 -309
rect 754 -392 764 -314
rect 876 -392 886 -314
rect 1006 -325 1011 -269
rect 1067 -325 1072 -269
rect 1006 -330 1072 -325
rect 754 -397 886 -392
rect 246 -484 316 -399
rect 792 -484 860 -397
rect 246 -500 860 -484
rect 247 -552 860 -500
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729243291
transform 1 0 1083 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729243291
transform 1 0 21 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729243291
transform 1 0 21 0 1 -329
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729243291
transform 1 0 1083 0 1 -329
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_BH5GQ5  sky130_fd_pr__pfet_01v8_BH5GQ5_1
timestamp 1729243291
transform 1 0 552 0 1 -329
box -552 -200 552 200
use sky130_fd_pr__pfet_01v8_BH5GQ5  sky130_fd_pr__pfet_01v8_BH5GQ5_2
timestamp 1729243291
transform 1 0 552 0 1 200
box -552 -200 552 200
<< labels >>
flabel viali 1228 -100 1228 -100 0 FreeSans 160 0 0 0 VDD
port 0 nsew
flabel via1 690 360 690 360 0 FreeSans 160 0 0 0 VIP
port 1 nsew
flabel via1 140 364 140 364 0 FreeSans 160 0 0 0 VIN
port 2 nsew
flabel via1 60 140 60 140 0 FreeSans 160 0 0 0 D6
port 3 nsew
flabel via2 62 -278 62 -278 0 FreeSans 160 0 0 0 D7
port 4 nsew
flabel metal1 262 32 262 32 0 FreeSans 1600 0 0 0 S
port 5 nsew
<< end >>
