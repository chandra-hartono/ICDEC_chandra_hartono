magic
tech sky130A
magscale 1 2
timestamp 1729156958
<< nwell >>
rect -39 247 977 3097
<< nsubdiff >>
rect -3 3027 57 3061
rect 881 3027 941 3061
rect -3 3001 31 3027
rect 907 3001 941 3027
rect -3 317 31 343
rect 907 317 941 343
rect -3 283 57 317
rect 881 283 941 317
<< nsubdiffcont >>
rect 57 3027 881 3061
rect -3 343 31 3001
rect 907 343 941 3001
rect 57 283 881 317
<< poly >>
rect 82 2961 174 2977
rect 82 2927 98 2961
rect 132 2927 174 2961
rect 82 2911 174 2927
rect 144 2904 174 2911
rect 746 2961 850 2976
rect 746 2927 790 2961
rect 824 2927 850 2961
rect 746 2896 850 2927
rect 81 2281 174 2297
rect 232 2292 432 2386
rect 81 2247 97 2281
rect 131 2247 174 2281
rect 81 2231 174 2247
rect 129 2224 174 2231
rect 748 2279 840 2296
rect 748 2245 790 2279
rect 824 2245 840 2279
rect 748 2223 840 2245
rect 83 1600 174 1616
rect 232 1610 690 1704
rect 83 1566 99 1600
rect 133 1566 174 1600
rect 83 1539 174 1566
rect 748 1599 836 1615
rect 748 1565 786 1599
rect 820 1565 836 1599
rect 748 1549 836 1565
rect 748 1543 835 1549
rect 78 917 174 933
rect 490 928 690 1024
rect 78 883 95 917
rect 129 883 174 917
rect 78 860 174 883
rect 748 917 841 933
rect 748 883 790 917
rect 824 883 841 917
rect 748 861 841 883
<< polycont >>
rect 98 2927 132 2961
rect 790 2927 824 2961
rect 97 2247 131 2281
rect 790 2245 824 2279
rect 99 1566 133 1600
rect 786 1565 820 1599
rect 95 883 129 917
rect 790 883 824 917
<< locali >>
rect -3 3027 57 3061
rect 881 3027 941 3061
rect -3 3001 31 3027
rect 907 3001 941 3027
rect 780 2961 834 2978
rect 82 2927 98 2961
rect 132 2927 148 2961
rect 780 2927 790 2961
rect 824 2927 834 2961
rect 98 2880 132 2927
rect 780 2918 834 2927
rect 788 2846 824 2918
rect 81 2247 97 2281
rect 131 2247 147 2281
rect 774 2274 790 2279
rect 90 2175 144 2247
rect 773 2245 790 2274
rect 824 2245 840 2279
rect 773 2183 831 2245
rect 706 2178 831 2183
rect 706 1821 824 2178
rect 83 1566 99 1600
rect 133 1566 149 1600
rect 94 1503 137 1566
rect 770 1565 786 1599
rect 820 1565 836 1599
rect 776 1486 835 1565
rect 79 883 95 917
rect 129 883 145 917
rect 774 883 790 917
rect 824 883 840 917
rect 84 814 137 883
rect 782 781 834 883
rect -3 317 31 343
rect 907 317 941 343
rect -3 283 57 317
rect 881 283 941 317
<< viali >>
rect 98 2927 132 2961
rect 790 2927 824 2961
rect 906 2920 907 2972
rect 907 2920 941 2972
rect 941 2920 942 2972
rect 97 2247 131 2281
rect 790 2245 824 2279
rect 99 1566 133 1600
rect 786 1565 820 1599
rect -4 874 -3 922
rect -3 874 30 922
rect 95 883 129 917
rect 790 883 824 917
<< metal1 >>
rect 780 2976 834 2978
rect 900 2976 948 2984
rect 780 2972 948 2976
rect 86 2961 226 2967
rect 86 2927 98 2961
rect 132 2927 226 2961
rect 86 2921 226 2927
rect 92 2880 138 2921
rect 180 2872 226 2921
rect 780 2961 906 2972
rect 780 2927 790 2961
rect 824 2927 906 2961
rect 780 2920 906 2927
rect 942 2920 948 2972
rect 780 2914 948 2920
rect 788 2871 826 2914
rect 900 2908 948 2914
rect 79 2492 89 2868
rect 141 2865 151 2868
rect 141 2554 218 2865
rect 141 2492 151 2554
rect 442 2431 478 2866
rect 691 2488 828 2871
rect 697 2431 738 2488
rect 442 2397 742 2431
rect 85 2281 143 2287
rect 85 2247 97 2281
rect 131 2252 143 2281
rect 131 2247 144 2252
rect 85 2241 144 2247
rect 90 2192 144 2241
rect 90 2175 219 2192
rect 94 2097 219 2175
rect 94 1838 182 2097
rect 234 1838 244 2097
rect 94 1809 219 1838
rect 87 1600 145 1606
rect 87 1566 99 1600
rect 133 1566 145 1600
rect 87 1560 145 1566
rect 187 1564 394 1601
rect 94 1512 137 1560
rect 187 1512 223 1564
rect 91 1128 228 1512
rect -10 922 36 934
rect 83 922 141 923
rect -10 874 -4 922
rect 30 917 141 922
rect 442 918 478 2397
rect 778 2279 836 2285
rect 778 2274 790 2279
rect 773 2245 790 2274
rect 824 2245 836 2279
rect 773 2239 836 2245
rect 773 2183 831 2239
rect 706 2178 831 2183
rect 706 1845 824 2178
rect 702 1821 824 1845
rect 702 1749 737 1821
rect 627 1713 737 1749
rect 774 1599 832 1605
rect 774 1565 786 1599
rect 820 1591 832 1599
rect 820 1565 835 1591
rect 774 1559 835 1565
rect 776 1511 835 1559
rect 696 1486 835 1511
rect 696 1468 831 1486
rect 683 1209 693 1468
rect 745 1209 831 1468
rect 696 1133 831 1209
rect 30 883 95 917
rect 129 883 141 917
rect 30 877 141 883
rect 186 916 218 918
rect 186 881 294 916
rect 390 882 479 918
rect 778 917 836 923
rect 778 883 790 917
rect 824 883 836 917
rect 30 874 138 877
rect -10 862 36 874
rect 84 821 137 874
rect 186 824 218 881
rect 186 821 220 824
rect 84 814 220 821
rect 91 459 220 814
rect 214 448 220 459
rect 442 448 478 882
rect 778 877 836 883
rect 782 826 834 877
rect 770 825 780 826
rect 703 584 780 825
rect 836 584 846 826
rect 703 461 825 584
<< via1 >>
rect 89 2492 141 2868
rect 182 1838 234 2097
rect 693 1209 745 1468
rect 780 584 836 826
<< metal2 >>
rect 89 2868 141 2878
rect 89 2482 141 2492
rect 97 2397 130 2482
rect 90 2364 150 2397
rect 90 2308 92 2364
rect 148 2308 150 2364
rect 90 1691 150 2308
rect 765 2306 774 2366
rect 834 2306 843 2366
rect 182 2097 234 2107
rect 182 1828 234 1838
rect 88 1682 150 1691
rect 148 1622 150 1682
rect 88 1620 150 1622
rect 183 1664 227 1828
rect 774 1680 834 2306
rect 183 1620 740 1664
rect 88 1004 148 1620
rect 696 1478 740 1620
rect 774 1624 776 1680
rect 832 1624 834 1680
rect 693 1468 745 1478
rect 693 1199 745 1209
rect 88 948 90 1004
rect 146 948 148 1004
rect 88 946 148 948
rect 774 1015 834 1624
rect 774 1006 838 1015
rect 774 946 778 1006
rect 90 939 146 946
rect 774 942 838 946
rect 778 937 838 942
rect 782 836 834 937
rect 780 826 836 836
rect 780 574 836 584
<< via2 >>
rect 92 2308 148 2364
rect 774 2306 834 2366
rect 88 1622 148 1682
rect 776 1624 832 1680
rect 90 948 146 1004
rect 778 946 838 1006
<< metal3 >>
rect 87 2366 153 2369
rect 769 2366 839 2371
rect 87 2364 774 2366
rect 87 2308 92 2364
rect 148 2308 774 2364
rect 87 2306 774 2308
rect 834 2306 839 2366
rect 87 2303 153 2306
rect 769 2301 839 2306
rect 83 1682 153 1687
rect 771 1682 837 1685
rect 83 1622 88 1682
rect 148 1680 837 1682
rect 148 1624 776 1680
rect 832 1624 837 1680
rect 148 1622 837 1624
rect 83 1617 153 1622
rect 771 1619 837 1622
rect 85 1006 151 1009
rect 773 1006 843 1011
rect 85 1004 778 1006
rect 85 948 90 1004
rect 146 948 778 1004
rect 85 946 778 948
rect 838 946 843 1006
rect 85 943 151 946
rect 773 941 843 946
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_8
timestamp 1729141747
transform 1 0 763 0 1 2680
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_9
timestamp 1729141747
transform 1 0 159 0 1 2680
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_10
timestamp 1729141747
transform 1 0 763 0 1 1998
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_11
timestamp 1729141747
transform 1 0 159 0 1 1998
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_12
timestamp 1729141747
transform 1 0 763 0 1 1318
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_13
timestamp 1729141747
transform 1 0 159 0 1 1318
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_14
timestamp 1729141747
transform 1 0 159 0 1 636
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_15
timestamp 1729141747
transform 1 0 763 0 1 636
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_4
timestamp 1729141747
transform 1 0 461 0 1 2680
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_5
timestamp 1729141747
transform 1 0 461 0 1 1998
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_6
timestamp 1729141747
transform 1 0 461 0 1 1318
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_7
timestamp 1729141747
transform 1 0 461 0 1 636
box -323 -300 323 300
<< labels >>
flabel metal1 868 2944 868 2944 0 FreeSans 160 0 0 0 VDD
port 0 nsew
flabel metal2 206 1722 206 1722 0 FreeSans 160 0 0 0 D1
port 1 nsew
flabel metal1 716 1734 716 1734 0 FreeSans 160 0 0 0 D2
port 2 nsew
flabel metal2 800 1722 800 1722 0 FreeSans 160 0 0 0 D5
port 3 nsew
<< end >>
