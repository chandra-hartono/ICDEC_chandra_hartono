magic
tech sky130A
magscale 1 2
timestamp 1729370620
<< psubdiff >>
rect -306 976 -246 1010
rect 1519 976 1579 1010
rect -306 933 -272 976
rect 1545 933 1579 976
rect -306 -191 -272 -103
rect 1545 -191 1579 -103
rect -306 -225 -246 -191
rect 1519 -225 1579 -191
<< psubdiffcont >>
rect -246 976 1519 1010
rect -306 -103 -272 933
rect 1545 -103 1579 933
rect -246 -225 1519 -191
<< poly >>
rect 56 326 1198 470
<< locali >>
rect -306 976 -246 1010
rect 1519 976 1579 1010
rect -306 933 -272 976
rect -306 -191 -272 -103
rect 1545 933 1579 976
rect 1545 -191 1579 -103
rect -306 -225 -246 -191
rect 1519 -225 1579 -191
<< viali >>
rect 914 976 1053 1010
rect 177 -225 333 -191
rect 177 -226 333 -225
<< metal1 >>
rect 902 1010 1065 1016
rect 902 976 914 1010
rect 1053 976 1065 1010
rect 902 970 1065 976
rect 928 932 1039 970
rect 594 848 1342 932
rect -188 744 -66 778
rect -188 676 -154 744
rect -100 694 -66 744
rect 594 694 678 848
rect 1258 778 1342 848
rect 1258 744 1460 778
rect 1258 694 1372 744
rect -100 575 46 694
rect -101 518 46 575
rect -101 276 -38 518
rect 246 462 281 540
rect 325 518 335 570
rect 387 518 397 570
rect 192 458 281 462
rect 189 434 281 458
rect 330 326 450 360
rect -206 50 -172 130
rect -120 100 46 276
rect 211 222 221 274
rect 273 222 283 274
rect 330 254 358 326
rect 586 100 686 694
rect 1224 572 1372 694
rect 1426 652 1460 744
rect 875 518 885 570
rect 937 518 947 570
rect 981 469 1023 544
rect 1224 518 1390 572
rect 981 435 1118 469
rect 981 434 1023 435
rect 843 326 946 360
rect 917 248 946 326
rect 988 226 998 278
rect 1050 226 1060 278
rect 1304 276 1390 518
rect 1226 100 1390 276
rect -118 50 -84 100
rect -206 16 -84 50
rect -39 -25 15 100
rect -38 -35 15 -25
rect 594 -35 680 100
rect 1356 50 1390 100
rect 1444 50 1478 102
rect 1356 16 1478 50
rect -38 -121 680 -35
rect 204 -185 307 -121
rect 165 -191 345 -185
rect 165 -226 177 -191
rect 333 -226 345 -191
rect 165 -232 345 -226
<< via1 >>
rect 335 518 387 570
rect 221 222 273 274
rect 885 518 937 570
rect 998 226 1050 278
<< metal2 >>
rect 335 570 387 580
rect 335 508 387 518
rect 885 570 937 580
rect 885 508 937 518
rect 344 414 380 508
rect 894 414 930 508
rect 344 413 930 414
rect 231 377 1041 413
rect 231 284 267 377
rect 1005 288 1041 377
rect 221 274 273 284
rect 221 212 273 222
rect 998 278 1050 288
rect 998 216 1050 226
use sky130_fd_pr__nfet_01v8_C77M8X  sky130_fd_pr__nfet_01v8_C77M8X_0
timestamp 1729360621
transform 1 0 636 0 1 397
box -636 -397 636 397
use sky130_fd_pr__nfet_01v8_UPT43B  sky130_fd_pr__nfet_01v8_UPT43B_0
timestamp 1729360787
transform 1 0 1417 0 -1 157
box -73 -157 73 157
use sky130_fd_pr__nfet_01v8_UPT43B  sky130_fd_pr__nfet_01v8_UPT43B_1
timestamp 1729360787
transform 1 0 -127 0 1 637
box -73 -157 73 157
use sky130_fd_pr__nfet_01v8_UPT43B  sky130_fd_pr__nfet_01v8_UPT43B_2
timestamp 1729360787
transform 1 0 1401 0 1 637
box -73 -157 73 157
use sky130_fd_pr__nfet_01v8_UPT43B  sky130_fd_pr__nfet_01v8_UPT43B_3
timestamp 1729360787
transform 1 0 -145 0 -1 157
box -73 -157 73 157
<< labels >>
flabel viali 948 996 948 996 0 FreeSans 320 0 0 0 GND
port 0 nsew
flabel metal1 262 516 262 516 0 FreeSans 320 0 0 0 D8
port 1 nsew
flabel via1 914 550 914 550 0 FreeSans 320 0 0 0 D9
port 2 nsew
<< end >>
