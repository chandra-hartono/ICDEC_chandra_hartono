magic
tech sky130A
magscale 1 2
timestamp 1729403493
<< metal1 >>
rect 940 2722 986 2724
rect 940 2668 1308 2722
rect 1254 2601 1308 2668
rect 1254 2547 1526 2601
rect 817 1744 3102 1798
rect 811 998 2291 1113
rect 3048 932 3102 1744
rect 2689 -52 2755 144
rect 1833 -304 1843 -247
rect 1904 -304 1914 -247
<< via1 >>
rect 1843 -304 1904 -247
<< metal2 >>
rect 2646 2872 2702 2874
rect 2636 2864 2702 2872
rect 3294 2866 3350 2872
rect 2636 2808 2646 2864
rect 2636 2780 2702 2808
rect 3291 2863 3353 2866
rect 3291 2807 3294 2863
rect 3350 2807 3353 2863
rect 3291 2756 3353 2807
rect 3291 2717 3357 2756
rect 817 1110 873 1116
rect 817 1040 873 1041
rect 1873 530 1950 2337
rect 820 517 1950 530
rect 820 436 1954 517
rect 3301 487 3357 2717
rect 820 422 1948 436
rect 3300 50 3357 487
rect 1847 -4 3357 50
rect 1847 -237 1901 -4
rect 3301 -5 3357 -4
rect 1843 -247 1904 -237
rect 1843 -314 1904 -304
rect 2735 -1379 2779 -754
rect 2735 -1388 2799 -1379
rect 2735 -1444 2743 -1388
rect 2735 -1453 2799 -1444
rect 2735 -1457 2779 -1453
<< via2 >>
rect 2646 2808 2702 2864
rect 3294 2807 3350 2863
rect 2743 -1444 2799 -1388
<< metal3 >>
rect 2636 2868 2712 2869
rect 2634 2866 2712 2868
rect 3289 2866 3355 2868
rect 2632 2864 3356 2866
rect 2632 2808 2646 2864
rect 2702 2863 3356 2864
rect 2702 2808 3294 2863
rect 2632 2807 3294 2808
rect 3350 2807 3356 2863
rect 2632 2804 3356 2807
rect 2634 2803 2712 2804
rect 2634 2790 2708 2803
rect 3289 2802 3355 2804
rect 2648 2355 3352 2415
rect 2738 -1386 2804 -1383
rect 3292 -1386 3352 2355
rect 2738 -1388 3352 -1386
rect 2738 -1444 2743 -1388
rect 2799 -1444 3352 -1388
rect 2738 -1446 3352 -1444
rect 2738 -1449 2804 -1446
use nmos34  nmos34_0
timestamp 1729223266
transform 1 0 2328 0 1 203
box -235 -98 869 1334
use nmos89  nmos89_0
timestamp 1729370620
transform 1 0 1738 0 1 -1036
box -306 -232 1579 1016
use pmos67  pmos67_0
timestamp 1729397135
transform -1 0 2740 0 1 2672
box -176 -694 1280 562
use pmoscs  pmoscs_0
timestamp 1729156958
transform 1 0 39 0 1 -247
box -39 247 977 3097
<< labels >>
flabel metal2 s 2698 3116 2698 3116 0 FreeSans 160 0 0 0 VIN
port 0 nsew
flabel metal2 s 1688 3114 1688 3116 0 FreeSans 160 0 0 0 VIP
port 1 nsew
flabel metal1 s 1210 2688 1210 2688 0 FreeSans 160 0 0 0 VDD
port 2 nsew
flabel metal1 s 2720 72 2720 72 0 FreeSans 160 0 0 0 GND
port 3 nsew
flabel metal3 s 2614 710 2614 710 0 FreeSans 160 0 0 0 RS
port 4 nsew
flabel metal3 s 3054 2390 3054 2390 0 FreeSans 160 0 0 0 OUT
port 5 nsew
<< end >>
